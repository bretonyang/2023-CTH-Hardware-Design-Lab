// StudentID StudentName

module exam1_A(a, b, c, d, sel, neg);
    input [2:0] a, b, c;
    input [1:0] sel;
    output neg;
    output [3:0] d;

    // add your design here

endmodule
