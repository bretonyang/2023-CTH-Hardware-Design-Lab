// StudentID StudentName

module exam1_B (clk, rst, Fn);
    input clk, rst;
    output [19:0] Fn;

    // add your design here
    
endmodule
