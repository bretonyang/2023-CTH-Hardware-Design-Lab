module clock_divider 
  #(parameter n = 25)
  (input clk, output clk_div);
  


endmodule