// 108123456 王小明
module exam2_A(clk, rst, en_btn, dir_btn, DIGIT, DISPLAY);
   input clk, rst, en_btn, dir_btn;
   output[3:0] DIGIT;
   output[6:0] DISPLAY;

   // add your design here
   
endmodule
